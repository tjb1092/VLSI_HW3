magic
tech scmos
timestamp 1538945983
<< ntransistor >>
rect 0 47 2 50
rect 32 47 34 50
rect 48 46 50 50
rect 64 47 66 50
rect 112 47 114 50
rect 80 41 82 45
rect 96 41 98 45
rect 112 33 114 37
rect 16 22 18 27
rect 32 22 34 27
rect 48 22 50 27
rect 64 22 66 27
rect 80 22 82 27
rect 0 9 2 14
rect 32 9 34 14
rect 48 9 50 14
rect 64 10 66 14
rect 80 10 82 14
<< ptransistor >>
rect 0 109 2 118
rect 32 107 34 117
rect 48 107 50 117
rect 64 107 66 117
rect 80 107 82 117
rect 16 94 18 103
rect 32 94 34 103
rect 48 94 50 103
rect 64 94 66 103
rect 80 94 82 103
rect 0 62 2 66
rect 48 75 50 82
rect 32 62 34 66
rect 80 70 82 77
rect 96 70 98 77
rect 112 70 114 77
rect 64 62 66 66
rect 112 62 114 66
<< ndiffusion >>
rect -1 47 0 50
rect 2 47 3 50
rect 31 47 32 50
rect 34 47 35 50
rect 47 46 48 50
rect 50 46 51 50
rect 63 47 64 50
rect 66 47 67 50
rect 111 47 112 50
rect 114 47 115 50
rect 79 41 80 45
rect 82 41 87 45
rect 91 41 96 45
rect 98 41 99 45
rect 111 33 112 37
rect 114 33 115 37
rect 15 23 16 27
rect 13 22 16 23
rect 18 23 19 27
rect 31 23 32 27
rect 18 22 21 23
rect 29 22 32 23
rect 34 23 39 27
rect 43 23 48 27
rect 34 22 48 23
rect 50 22 64 27
rect 66 23 71 27
rect 75 23 80 27
rect 66 22 80 23
rect 82 23 83 27
rect 82 22 85 23
rect -1 10 0 14
rect -3 9 0 10
rect 2 10 3 14
rect 2 9 5 10
rect 31 10 32 14
rect 29 9 32 10
rect 34 10 39 14
rect 43 10 48 14
rect 34 9 48 10
rect 50 10 51 14
rect 63 10 64 14
rect 66 10 71 14
rect 75 10 80 14
rect 82 10 83 14
rect 50 9 53 10
<< pdiffusion >>
rect -3 113 0 118
rect -1 109 0 113
rect 2 116 7 118
rect 2 112 3 116
rect 2 109 7 112
rect 29 112 32 117
rect 31 108 32 112
rect 27 107 32 108
rect 34 115 48 117
rect 34 111 39 115
rect 43 111 48 115
rect 34 107 48 111
rect 50 107 64 117
rect 66 115 80 117
rect 66 111 71 115
rect 75 111 80 115
rect 66 107 80 111
rect 82 112 85 117
rect 82 108 83 112
rect 82 107 87 108
rect 13 98 16 103
rect 15 94 16 98
rect 18 98 32 103
rect 18 94 23 98
rect 27 94 32 98
rect 34 98 48 103
rect 34 94 39 98
rect 43 94 48 98
rect 50 101 64 103
rect 50 97 55 101
rect 59 97 64 101
rect 50 94 64 97
rect 66 98 80 103
rect 66 94 71 98
rect 75 94 80 98
rect 82 98 85 103
rect 82 94 83 98
rect -1 62 0 66
rect 2 62 3 66
rect 45 79 48 82
rect 47 75 48 79
rect 50 79 53 82
rect 50 75 51 79
rect 31 62 32 66
rect 34 62 35 66
rect 77 74 80 77
rect 79 70 80 74
rect 82 70 96 77
rect 98 74 112 77
rect 98 70 105 74
rect 109 70 112 74
rect 114 73 115 77
rect 114 70 119 73
rect 63 62 64 66
rect 66 62 67 66
rect 111 62 112 66
rect 114 62 115 66
<< ndcontact >>
rect -5 46 -1 50
rect 3 46 7 50
rect 27 46 31 50
rect 35 46 39 50
rect 43 46 47 50
rect 51 46 55 50
rect 59 46 63 50
rect 67 46 71 50
rect 107 46 111 50
rect 75 41 79 45
rect 87 41 91 45
rect 99 41 103 45
rect 115 46 119 50
rect 107 33 111 37
rect 115 33 119 37
rect 11 23 15 27
rect 19 23 23 27
rect 27 23 31 27
rect 39 23 43 27
rect 71 23 75 27
rect 83 23 87 27
rect -5 10 -1 14
rect 3 10 7 14
rect 27 10 31 14
rect 39 10 43 14
rect 51 10 55 14
rect 59 10 63 14
rect 71 10 75 14
rect 83 10 87 14
<< pdcontact >>
rect -5 109 -1 113
rect 3 112 7 116
rect 27 108 31 112
rect 39 111 43 115
rect 71 111 75 115
rect 83 108 87 112
rect 11 94 15 98
rect 23 94 27 98
rect 39 94 43 98
rect 55 97 59 101
rect 71 94 75 98
rect 83 94 87 98
rect -5 62 -1 66
rect 3 62 7 66
rect 43 75 47 79
rect 51 75 55 79
rect 27 62 31 66
rect 35 62 39 66
rect 75 70 79 74
rect 105 70 109 74
rect 115 73 119 77
rect 59 62 63 66
rect 67 62 71 66
rect 107 62 111 66
rect 115 62 119 66
<< polysilicon >>
rect 0 118 2 128
rect 0 66 2 109
rect 16 103 18 121
rect 32 117 34 134
rect 48 117 50 121
rect 64 117 66 134
rect 80 117 82 121
rect 32 103 34 107
rect 48 103 50 107
rect 64 103 66 107
rect 80 103 82 107
rect 0 50 2 62
rect 16 58 18 94
rect 32 66 34 94
rect 48 82 50 94
rect 17 54 18 58
rect 0 14 2 47
rect 16 27 18 54
rect 32 50 34 62
rect 48 61 50 75
rect 64 66 66 94
rect 80 77 82 94
rect 96 77 98 87
rect 112 77 114 87
rect 49 57 50 61
rect 48 50 50 57
rect 64 50 66 62
rect 80 58 82 70
rect 81 54 82 58
rect 32 27 34 47
rect 48 27 50 46
rect 64 27 66 47
rect 80 45 82 54
rect 96 58 98 70
rect 112 66 114 70
rect 96 54 97 58
rect 96 45 98 54
rect 112 50 114 62
rect 80 27 82 41
rect 96 34 98 41
rect 112 37 114 47
rect 0 7 2 9
rect 16 7 18 22
rect 32 14 34 22
rect 48 14 50 22
rect 64 14 66 22
rect 80 14 82 22
rect 32 7 34 9
rect 48 7 50 9
rect 64 7 66 10
rect 80 7 82 10
rect 112 0 114 33
<< polycontact >>
rect 31 134 35 138
rect 63 134 67 138
rect -1 128 3 132
rect 13 54 17 58
rect 45 57 49 61
rect 77 54 81 58
rect 97 54 101 58
rect 111 -4 115 0
<< metal1 >>
rect -16 128 -11 131
rect 3 128 129 131
rect -16 121 129 125
rect -13 72 -10 121
rect 4 116 43 118
rect 7 115 43 116
rect -5 98 -2 109
rect 55 101 58 121
rect 71 115 74 121
rect -3 97 -2 98
rect -3 94 11 97
rect 40 91 43 94
rect 71 91 74 94
rect 40 88 74 91
rect 44 82 118 85
rect 44 79 47 82
rect 52 72 55 75
rect 115 77 118 82
rect -13 70 75 72
rect -13 69 79 70
rect -4 66 -1 69
rect 27 66 30 69
rect 60 66 63 69
rect 122 66 125 121
rect 4 57 7 62
rect 36 60 39 62
rect 4 54 13 57
rect 36 57 45 60
rect 68 57 71 62
rect 119 63 125 66
rect 4 50 7 54
rect 36 50 39 57
rect 68 54 77 57
rect 107 57 110 62
rect 101 54 110 57
rect 68 50 71 54
rect -5 43 -2 46
rect 27 43 30 46
rect -5 40 30 43
rect 107 50 110 54
rect 119 46 129 49
rect -5 14 -2 40
rect 59 37 62 46
rect 76 37 79 41
rect 126 43 129 46
rect 103 41 129 43
rect 99 40 129 41
rect 11 34 42 37
rect 59 34 93 37
rect 11 27 14 34
rect 39 27 42 34
rect 75 23 80 26
rect 20 13 23 23
rect 77 20 80 23
rect 40 17 74 20
rect 77 18 87 20
rect 77 17 83 18
rect 40 14 43 17
rect 71 14 74 17
rect 7 10 27 13
rect -5 7 -2 10
rect 52 7 55 10
rect 59 7 62 10
rect 90 7 93 34
rect 126 7 129 40
rect -16 3 129 7
rect -16 -3 111 0
rect 115 -3 129 0
<< m2contact >>
rect -11 128 -7 132
rect 27 104 31 108
rect 83 104 87 108
rect -7 94 -3 98
rect 23 90 27 94
rect 83 90 87 94
rect 101 70 105 74
rect 43 50 47 54
rect 51 42 55 46
rect 91 40 95 44
rect 7 33 11 37
rect 27 27 31 31
rect 83 27 87 31
rect 27 14 31 18
rect 83 14 87 18
rect 103 33 107 37
rect 119 33 123 37
rect 119 -10 123 -6
<< metal2 >>
rect -10 37 -7 128
rect 31 105 83 108
rect 27 91 83 94
rect 101 69 104 70
rect 92 66 104 69
rect 92 53 95 66
rect 47 50 122 53
rect 52 40 55 42
rect 52 37 107 40
rect -10 34 7 37
rect 119 37 122 50
rect 31 27 83 30
rect 31 14 83 17
rect 119 -6 122 33
<< labels >>
rlabel polysilicon 64 7 66 10 1 b
rlabel polysilicon 80 7 82 10 1 bbar
rlabel polysilicon 96 34 98 37 1 minbar
rlabel polysilicon 112 30 114 33 1 min
rlabel polysilicon 16 7 18 10 1 pinbar
rlabel metal1 -5 121 -3 123 1 vdd
rlabel metal1 -16 128 -14 130 3 pout
rlabel metal1 -3 3 -1 5 1 gnd
rlabel metal2 119 -6 121 -4 1 fout
rlabel polysilicon 48 7 50 9 1 abar
rlabel polysilicon 32 131 34 133 1 a
rlabel polysilicon 0 125 2 127 1 pin
<< end >>
