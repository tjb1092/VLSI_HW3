magic
tech scmos
timestamp 1538870037
<< ntransistor >>
rect -6 12 -4 16
rect 10 12 12 16
rect 58 20 60 23
rect 74 12 76 15
rect 122 20 124 24
rect 138 20 140 24
rect 154 20 156 24
rect 122 12 124 16
rect 138 12 140 16
rect 26 4 28 8
rect 42 4 44 8
rect 58 4 60 8
rect 74 4 76 8
rect 90 4 92 8
rect 106 4 108 8
rect 122 4 124 8
rect 138 4 140 8
rect 154 4 156 8
rect 170 4 172 8
rect 186 4 188 8
rect 202 4 204 8
<< ptransistor >>
rect 122 65 124 69
rect 138 65 140 69
rect -6 52 -4 56
rect 10 52 12 56
rect 26 52 28 56
rect 42 52 44 56
rect 58 52 60 56
rect 74 52 76 56
rect 90 52 92 56
rect 106 52 108 56
rect 122 52 124 56
rect 138 52 140 56
rect 154 52 156 56
rect 170 52 172 56
rect 58 36 60 40
rect 74 36 76 40
rect 122 38 124 42
rect 138 36 140 40
rect 154 36 156 40
rect 186 36 188 40
rect 202 36 204 40
<< ndiffusion >>
rect -7 12 -6 16
rect -4 12 10 16
rect 12 12 13 16
rect 57 20 58 23
rect 60 20 61 23
rect 73 12 74 15
rect 76 12 77 15
rect 121 20 122 24
rect 124 20 125 24
rect 137 20 138 24
rect 140 20 141 24
rect 153 20 154 24
rect 156 20 157 24
rect 121 12 122 16
rect 124 12 127 16
rect 131 12 138 16
rect 140 12 141 16
rect 25 4 26 8
rect 28 4 42 8
rect 44 4 45 8
rect 57 4 58 8
rect 60 4 74 8
rect 76 4 77 8
rect 89 4 90 8
rect 92 4 97 8
rect 101 4 106 8
rect 108 4 109 8
rect 121 4 122 8
rect 124 4 125 8
rect 137 4 138 8
rect 140 4 154 8
rect 156 4 157 8
rect 169 4 170 8
rect 172 4 173 8
rect 185 4 186 8
rect 188 4 202 8
rect 204 4 205 8
<< pdiffusion >>
rect 121 65 122 69
rect 124 65 125 69
rect 137 65 138 69
rect 140 65 141 69
rect -7 52 -6 56
rect -4 52 -3 56
rect 9 52 10 56
rect 12 52 13 56
rect 25 52 26 56
rect 28 52 29 56
rect 41 52 42 56
rect 44 52 45 56
rect 57 52 58 56
rect 60 52 61 56
rect 73 52 74 56
rect 76 52 77 56
rect 89 52 90 56
rect 92 52 93 56
rect 105 52 106 56
rect 108 52 109 56
rect 121 52 122 56
rect 124 52 125 56
rect 137 52 138 56
rect 140 52 141 56
rect 153 52 154 56
rect 156 52 157 56
rect 169 52 170 56
rect 172 52 173 56
rect 57 36 58 40
rect 60 36 61 40
rect 73 36 74 40
rect 76 36 77 40
rect 117 38 122 42
rect 124 38 125 42
rect 137 36 138 40
rect 140 36 141 40
rect 153 36 154 40
rect 156 36 157 40
rect 185 36 186 40
rect 188 36 189 40
rect 201 36 202 40
rect 204 36 205 40
<< ndcontact >>
rect -11 12 -7 16
rect 13 12 17 16
rect 53 20 57 24
rect 61 20 65 24
rect 69 12 73 16
rect 77 12 81 16
rect 117 20 121 24
rect 125 20 129 24
rect 133 20 137 24
rect 141 20 145 24
rect 149 20 153 24
rect 157 20 161 24
rect 117 12 121 16
rect 127 12 131 16
rect 141 12 145 16
rect 21 4 25 8
rect 45 4 49 8
rect 53 4 57 8
rect 77 4 81 8
rect 85 4 89 8
rect 97 4 101 8
rect 109 4 113 8
rect 117 4 121 8
rect 125 4 129 8
rect 133 4 137 8
rect 157 4 161 8
rect 165 4 169 8
rect 173 4 177 8
rect 181 4 185 8
rect 205 4 209 8
<< pdcontact >>
rect 117 65 121 69
rect 125 65 129 69
rect 133 65 137 69
rect 141 65 145 69
rect -11 52 -7 56
rect -3 52 1 56
rect 5 52 9 56
rect 13 52 17 56
rect 21 52 25 56
rect 29 52 33 56
rect 37 52 41 56
rect 45 52 49 56
rect 53 52 57 56
rect 61 52 65 56
rect 69 52 73 56
rect 77 52 81 56
rect 85 52 89 56
rect 93 52 97 56
rect 101 52 105 56
rect 109 52 113 56
rect 117 52 121 56
rect 125 52 129 56
rect 133 52 137 56
rect 141 52 145 56
rect 149 52 153 56
rect 157 52 161 56
rect 165 52 169 56
rect 173 52 177 56
rect 53 36 57 40
rect 61 36 65 40
rect 69 36 73 40
rect 77 36 81 40
rect 113 38 117 42
rect 125 38 129 42
rect 133 36 137 40
rect 141 36 145 40
rect 149 36 153 40
rect 157 36 161 40
rect 181 36 185 40
rect 189 36 193 40
rect 197 36 201 40
rect 205 36 209 40
<< polysilicon >>
rect -6 56 -4 59
rect 10 56 12 58
rect 26 56 28 58
rect 42 56 44 58
rect 58 56 60 83
rect 122 69 124 89
rect 138 69 140 89
rect 74 56 76 58
rect 90 56 92 58
rect 106 56 108 58
rect 122 56 124 65
rect 138 56 140 65
rect 154 56 156 58
rect 170 56 172 58
rect -6 32 -4 52
rect 10 32 12 52
rect -6 28 -5 32
rect 10 28 11 32
rect -6 16 -4 28
rect 10 16 12 28
rect 26 24 28 52
rect 42 35 44 52
rect 58 40 60 52
rect 74 40 76 52
rect 42 31 43 35
rect -6 -1 -4 12
rect 10 -2 12 12
rect 26 8 28 20
rect 42 8 44 31
rect 58 23 60 36
rect 74 27 76 36
rect 90 35 92 52
rect 90 31 91 35
rect 74 23 75 27
rect 58 8 60 20
rect 74 15 76 23
rect 74 8 76 12
rect 90 8 92 31
rect 106 27 108 52
rect 122 42 124 52
rect 138 40 140 52
rect 154 40 156 52
rect 106 23 107 27
rect 122 24 124 38
rect 138 24 140 36
rect 154 24 156 36
rect 170 35 172 52
rect 186 40 188 58
rect 202 40 204 58
rect 171 31 172 35
rect 106 8 108 23
rect 122 16 124 20
rect 138 16 140 20
rect 122 8 124 12
rect 138 8 140 12
rect 154 8 156 20
rect 170 8 172 31
rect 186 24 188 36
rect 202 24 204 36
rect 187 20 188 24
rect 203 20 204 24
rect 186 8 188 20
rect 202 8 204 20
rect 26 -2 28 4
rect 42 -2 44 4
rect 58 -2 60 4
rect 74 -2 76 4
rect 90 -2 92 4
rect 106 -2 108 4
rect 122 -2 124 4
rect 138 -2 140 4
rect 154 -17 156 4
rect 170 -2 172 4
rect 186 -2 188 4
rect 202 -2 204 4
<< polycontact >>
rect 121 89 125 93
rect 137 89 141 93
rect 57 83 61 87
rect -5 28 -1 32
rect 11 28 15 32
rect 43 31 47 35
rect 26 20 30 24
rect 91 31 95 35
rect 75 23 79 27
rect 107 23 111 27
rect 167 31 171 35
rect 183 20 187 24
rect 199 20 203 24
rect 153 -21 157 -17
<< metal1 >>
rect -17 83 -10 86
rect 61 83 214 86
rect -17 76 214 80
rect -10 59 8 62
rect -10 56 -7 59
rect 5 56 8 59
rect 13 56 16 76
rect 22 59 40 62
rect 54 59 72 62
rect 22 56 25 59
rect 37 56 40 59
rect 54 56 57 59
rect 69 56 72 59
rect 78 56 81 76
rect 126 69 129 76
rect 129 65 133 68
rect 145 65 160 68
rect 133 62 136 65
rect 94 59 120 62
rect 94 56 97 59
rect 117 56 120 59
rect 126 59 144 62
rect 126 56 129 59
rect 141 56 144 59
rect 157 56 160 65
rect 165 56 168 76
rect -11 16 -8 52
rect -2 49 1 52
rect 13 49 16 52
rect -2 46 16 49
rect 21 43 24 52
rect 30 49 33 52
rect 46 49 49 52
rect 62 49 65 52
rect 78 49 81 52
rect 30 46 81 49
rect 2 40 24 43
rect 2 31 5 40
rect 62 40 65 46
rect 78 40 81 46
rect -1 28 5 31
rect 37 31 40 39
rect 145 53 149 56
rect 85 49 88 52
rect 101 49 104 52
rect 85 46 104 49
rect 110 49 113 52
rect 133 49 136 52
rect 110 46 136 49
rect 53 34 56 36
rect 47 31 56 34
rect 15 28 40 31
rect 2 22 5 28
rect 2 19 23 22
rect 13 -10 16 12
rect 20 8 23 19
rect 37 14 40 28
rect 53 24 56 31
rect 37 11 56 14
rect 53 8 56 11
rect 20 4 21 8
rect 46 1 49 4
rect 62 1 65 20
rect 69 16 72 36
rect 85 26 88 46
rect 142 40 145 52
rect 157 46 160 52
rect 157 43 177 46
rect 114 27 117 38
rect 145 37 149 40
rect 79 23 88 26
rect 111 24 120 27
rect 85 15 88 23
rect 133 24 136 36
rect 158 34 161 36
rect 158 31 167 34
rect 158 24 161 31
rect 145 20 149 23
rect 174 23 177 43
rect 190 43 209 46
rect 190 40 193 43
rect 206 40 209 43
rect 181 33 184 36
rect 197 33 200 36
rect 181 30 200 33
rect 174 20 183 23
rect 206 24 209 36
rect 190 20 199 23
rect 206 20 207 24
rect 141 16 144 20
rect 164 17 177 20
rect 85 12 117 15
rect 164 14 167 17
rect 190 14 193 20
rect 46 -2 65 1
rect 77 8 80 12
rect 85 8 88 12
rect 141 8 144 12
rect 158 11 167 14
rect 174 11 193 14
rect 158 8 161 11
rect 174 8 177 11
rect 206 8 209 20
rect 113 4 117 7
rect 137 5 144 8
rect 54 -10 57 -2
rect 77 -10 80 4
rect 117 -10 120 4
rect 126 -3 129 4
rect 134 -10 137 4
rect 181 -10 184 4
rect -17 -14 214 -10
rect -17 -20 153 -17
rect 157 -20 214 -17
<< m2contact >>
rect -10 83 -6 87
rect -10 62 -6 66
rect 50 59 54 63
rect 97 72 101 76
rect 117 69 121 73
rect 37 39 41 43
rect 177 52 181 56
rect 30 20 34 24
rect 65 27 69 31
rect 121 38 125 42
rect 95 31 99 35
rect 129 31 133 35
rect 125 24 129 28
rect 141 24 145 28
rect 190 23 194 27
rect 207 20 211 24
rect 131 12 135 16
rect 97 0 101 4
rect 126 -7 130 -3
rect 165 0 169 4
rect 210 -27 214 -23
<< metal2 >>
rect 57 84 61 87
rect -10 66 -7 83
rect 50 43 53 59
rect 41 40 53 43
rect 98 45 101 72
rect 121 70 180 73
rect 177 56 180 70
rect 98 42 124 45
rect 99 32 129 35
rect 47 27 65 30
rect 47 24 50 27
rect 129 24 141 27
rect 177 27 180 52
rect 177 24 190 27
rect 26 21 30 24
rect 34 21 50 24
rect 131 3 134 12
rect 101 0 134 3
rect 165 -3 168 0
rect 130 -6 168 -3
rect 153 -20 157 -17
rect 211 -23 214 23
<< labels >>
rlabel polysilicon 26 -1 28 2 1 sbar
rlabel polysilicon 42 -1 44 2 1 pinb
rlabel polysilicon 58 -1 60 2 1 pin
rlabel polysilicon 74 -1 76 2 1 s
rlabel polysilicon 90 -1 92 2 1 bbar
rlabel polysilicon 106 -1 108 2 1 abar
rlabel polysilicon 122 -2 124 0 1 a
rlabel polysilicon 138 -2 140 0 1 b
rlabel polysilicon 154 -2 156 0 1 min
rlabel polysilicon 170 -2 172 1 1 minbar
rlabel polysilicon 186 -2 188 1 1 f3
rlabel polysilicon 202 -2 204 1 1 f4
rlabel polysilicon 10 -1 12 3 1 f1
rlabel polysilicon -6 0 -4 4 1 f2
<< end >>
