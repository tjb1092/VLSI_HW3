magic
tech scmos
timestamp 1539028648
<< ntransistor >>
rect 0 47 2 50
rect 32 45 34 50
rect 64 45 66 50
rect 48 31 50 35
rect 96 47 98 50
rect 80 31 82 35
rect 96 31 98 35
rect 112 31 114 35
rect 16 22 18 27
rect 32 22 34 27
rect 48 22 50 27
rect 64 22 66 27
rect 80 22 82 27
rect 0 9 2 14
rect 32 9 34 14
rect 48 9 50 14
rect 64 9 66 14
rect 80 9 82 14
<< ptransistor >>
rect 0 100 2 109
rect 32 101 34 110
rect 48 101 50 110
rect 64 101 66 110
rect 80 101 82 110
rect 16 86 18 95
rect 32 86 34 95
rect 48 86 50 95
rect 64 86 66 95
rect 80 86 82 95
rect 0 62 2 66
rect 48 74 50 82
rect 32 62 34 69
rect 80 70 82 78
rect 96 70 98 78
rect 112 70 114 78
rect 64 62 66 69
rect 96 62 98 66
<< ndiffusion >>
rect -1 47 0 50
rect 2 47 3 50
rect 31 46 32 50
rect 29 45 32 46
rect 34 46 35 50
rect 34 45 37 46
rect 63 46 64 50
rect 61 45 64 46
rect 66 46 67 50
rect 66 45 69 46
rect 47 31 48 35
rect 50 31 51 35
rect 95 47 96 50
rect 98 47 99 50
rect 79 31 80 35
rect 82 31 91 35
rect 95 31 96 35
rect 98 31 105 35
rect 109 31 112 35
rect 114 31 115 35
rect 15 23 16 27
rect 13 22 16 23
rect 18 23 19 27
rect 31 23 32 27
rect 18 22 21 23
rect 29 22 32 23
rect 34 23 36 27
rect 40 23 48 27
rect 34 22 48 23
rect 50 22 64 27
rect 66 23 71 27
rect 75 23 80 27
rect 66 22 80 23
rect 82 23 83 27
rect 82 22 85 23
rect -1 10 0 14
rect -3 9 0 10
rect 2 10 3 14
rect 31 10 32 14
rect 2 9 5 10
rect 29 9 32 10
rect 34 10 39 14
rect 43 10 48 14
rect 34 9 48 10
rect 50 10 51 14
rect 63 10 64 14
rect 50 9 53 10
rect 60 9 64 10
rect 66 10 71 14
rect 75 10 80 14
rect 66 9 80 10
rect 82 10 83 14
rect 82 9 85 10
<< pdiffusion >>
rect -3 104 0 109
rect -1 100 0 104
rect 2 106 3 109
rect 2 100 5 106
rect 29 105 32 110
rect 31 101 32 105
rect 34 107 35 110
rect 39 107 48 110
rect 34 101 48 107
rect 50 101 64 110
rect 66 107 71 110
rect 75 107 80 110
rect 66 101 80 107
rect 82 105 85 110
rect 82 101 83 105
rect 15 91 16 95
rect 13 86 16 91
rect 18 90 32 95
rect 18 86 27 90
rect 31 86 32 90
rect 34 90 48 95
rect 34 86 43 90
rect 47 86 48 90
rect 50 93 55 95
rect 59 93 64 95
rect 50 86 64 93
rect 66 90 80 95
rect 66 86 67 90
rect 71 86 80 90
rect 82 90 85 95
rect 82 86 83 90
rect -1 62 0 66
rect 2 62 3 66
rect 45 79 48 82
rect 47 75 48 79
rect 45 74 48 75
rect 50 80 53 82
rect 50 76 51 80
rect 50 74 53 76
rect 29 66 32 69
rect 31 62 32 66
rect 34 66 37 69
rect 34 62 35 66
rect 77 74 80 78
rect 79 70 80 74
rect 82 70 96 78
rect 98 74 112 78
rect 98 70 101 74
rect 105 70 112 74
rect 114 74 115 78
rect 114 70 119 74
rect 61 66 64 69
rect 63 62 64 66
rect 66 66 69 69
rect 66 62 67 66
rect 95 62 96 66
rect 98 62 99 66
<< ndcontact >>
rect -5 46 -1 50
rect 3 46 7 50
rect 27 46 31 50
rect 35 46 39 50
rect 59 46 63 50
rect 67 46 71 50
rect 43 31 47 35
rect 51 31 55 35
rect 91 46 95 50
rect 99 46 103 50
rect 75 31 79 35
rect 91 31 95 35
rect 105 31 109 35
rect 115 31 119 35
rect 11 23 15 27
rect 19 23 23 27
rect 27 23 31 27
rect 36 23 40 27
rect 71 23 75 27
rect 83 23 87 27
rect -5 10 -1 14
rect 3 10 7 14
rect 27 10 31 14
rect 39 10 43 14
rect 51 10 55 14
rect 59 10 63 14
rect 71 10 75 14
rect 83 10 87 14
<< pdcontact >>
rect -5 100 -1 104
rect 3 106 7 110
rect 27 101 31 105
rect 35 107 39 111
rect 71 107 75 111
rect 83 101 87 105
rect 11 91 15 95
rect 27 86 31 90
rect 43 86 47 90
rect 55 93 59 97
rect 67 86 71 90
rect 83 86 87 90
rect -5 62 -1 66
rect 3 62 7 66
rect 43 75 47 79
rect 51 76 55 80
rect 27 62 31 66
rect 35 62 39 66
rect 75 70 79 74
rect 101 70 105 74
rect 115 74 119 78
rect 59 62 63 66
rect 67 62 71 66
rect 91 62 95 66
rect 99 62 103 66
<< polysilicon >>
rect 0 109 2 121
rect 32 110 34 127
rect 48 110 50 113
rect 64 110 66 127
rect 80 110 82 113
rect 0 66 2 100
rect 16 95 18 98
rect 32 95 34 101
rect 48 95 50 101
rect 64 95 66 101
rect 80 95 82 101
rect 0 50 2 62
rect 16 58 18 86
rect 32 69 34 86
rect 48 82 50 86
rect 17 54 18 58
rect 0 14 2 47
rect 16 27 18 54
rect 32 50 34 62
rect 48 58 50 74
rect 64 69 66 86
rect 80 78 82 86
rect 96 78 98 80
rect 112 78 114 80
rect 49 54 50 58
rect 32 27 34 45
rect 48 35 50 54
rect 64 50 66 62
rect 80 58 82 70
rect 96 66 98 70
rect 81 54 82 58
rect 48 27 50 31
rect 64 27 66 45
rect 80 35 82 54
rect 96 50 98 62
rect 112 58 114 70
rect 113 54 114 58
rect 96 35 98 47
rect 112 35 114 54
rect 80 27 82 31
rect 16 19 18 22
rect 32 14 34 22
rect 48 14 50 22
rect 64 14 66 22
rect 80 14 82 22
rect 0 7 2 9
rect 32 7 34 9
rect 48 7 50 9
rect 64 7 66 9
rect 80 7 82 9
rect 96 0 98 31
rect 112 28 114 31
<< polycontact >>
rect 31 127 35 131
rect 63 127 67 131
rect -1 121 3 125
rect 13 54 17 58
rect 45 54 49 58
rect 77 54 81 58
rect 109 54 113 58
rect 95 -4 99 0
<< metal1 >>
rect -16 121 -11 124
rect 3 121 123 124
rect -16 114 123 118
rect -13 72 -10 114
rect 3 110 35 111
rect 7 108 35 110
rect -5 95 -2 100
rect 55 97 58 114
rect 71 111 74 114
rect -1 91 11 94
rect 47 86 67 89
rect 55 78 119 80
rect 55 77 115 78
rect 43 72 46 75
rect -13 70 75 72
rect -13 69 79 70
rect -4 66 -1 69
rect 27 66 30 69
rect 60 66 63 69
rect 76 66 79 69
rect 76 63 91 66
rect 4 57 7 62
rect 4 54 13 57
rect 36 57 39 62
rect 36 54 45 57
rect 68 57 71 62
rect 68 54 77 57
rect 100 57 103 62
rect 100 54 109 57
rect 4 50 7 54
rect 36 50 39 54
rect 68 50 71 54
rect 100 50 103 54
rect -5 43 -2 46
rect 27 43 30 46
rect -5 40 30 43
rect 60 43 63 46
rect 91 43 94 46
rect 60 40 94 43
rect -5 14 -2 40
rect 11 34 39 37
rect 11 27 14 34
rect 36 27 39 34
rect 55 33 58 34
rect 91 35 94 40
rect 62 33 75 34
rect 55 31 75 33
rect 75 23 80 26
rect 20 13 23 23
rect 77 20 80 23
rect 40 17 74 20
rect 77 18 87 20
rect 77 17 83 18
rect 40 14 43 17
rect 71 14 74 17
rect 7 10 27 13
rect -5 7 -2 10
rect 52 7 55 10
rect 59 7 62 10
rect 91 7 94 31
rect -16 3 123 7
rect -16 -3 95 0
rect 99 -3 123 0
<< m2contact >>
rect -11 121 -7 125
rect 27 97 31 101
rect 83 97 87 101
rect -5 91 -1 95
rect 27 90 31 94
rect 83 90 87 94
rect 105 70 109 74
rect 7 33 11 37
rect 27 27 31 31
rect 43 35 47 39
rect 58 33 62 37
rect 101 31 105 35
rect 119 31 123 35
rect 83 27 87 31
rect 27 14 31 18
rect 83 14 87 18
rect 119 -10 123 -6
<< metal2 >>
rect -10 95 -7 121
rect 31 98 83 101
rect -10 91 -5 95
rect -10 37 -7 91
rect 31 90 83 93
rect 106 67 109 70
rect 106 64 122 67
rect 119 44 122 64
rect 44 41 122 44
rect 44 39 47 41
rect -10 34 7 37
rect 58 37 105 38
rect 62 35 105 37
rect 119 35 122 41
rect 31 27 83 30
rect 31 14 83 17
rect 119 -6 122 31
<< labels >>
rlabel metal1 -3 3 -1 5 1 gnd
rlabel metal2 119 -6 121 -4 1 fout
rlabel polysilicon 48 7 50 9 1 abar
rlabel metal1 -15 121 -13 123 3 pout
rlabel polysilicon 0 118 2 120 1 pin
rlabel polysilicon 32 124 34 126 1 a
rlabel polysilicon 96 0 98 2 1 min
rlabel polysilicon 112 38 114 40 1 minbar
rlabel polysilicon 64 124 66 126 1 b
rlabel metal1 -15 114 -13 116 3 vdd
rlabel polysilicon 16 19 18 22 1 pinbar
rlabel polysilicon 80 7 82 9 1 bbar
<< end >>
