* SPICE3 file created from P3_take2.ext - technology: scmos

***************************************************
.include /home/baileytj/MOSFET_Models/IntroToVLSI/model_t36s.sp

.option scale=0.3u
.param vdd=5V

***************************************************
* Voltage Sources

vdd vdd 0 vdd
Vpin pin 0 PWL(0 0V 100n 0V 100.1n 0V 200n 0V 200.1n 0V 300n 0V 300.1n 0V 400n 0V 400.1n 0V 
+ 500n 0V 500.1n 0V 600n 0V 600.1n 0V 700n 0V 700.1n 0V 800n 0V 800.1n 5V 900n 5V 900.1n 5V 
+ 1000n 5V 1000.1n 5V 1100n 5V 1100.1n 5V 1200n 5V 1200.1n 5V 1300n 5V 1300.1n 5V 1400n 5V 1400.1n 5V 
+ 1500n 5V 1500.1n 5V 1600n 5V 1600.1n 5V 1700n 5V 1700.1n 0V)
A
Vmin min 0 PWL(0 0V 100n 0V 100.1n 0V 200n 0V 200.1n 0V 300n 0V 300.1n 0V 400n 0V 400.1n 0V 
+ 500n 0V 500.1n 0V 600n 0V 600.1n 0V 700n 0V 700.1n 0V 800n 0V 800.1n 5V 900n 5V 900.1n 5V 
+ 1000n 5V 1000.1n 5V 1100n 5V 1100.1n 5V 1200n 5V 1200.1n 5V 1300n 5V 1300.1n 5V 1400n 5V 1400.1n 5V 
+ 1500n 5V 1500.1n 5V 1600n 5V 1600.1n 5V 1700n 5V 1700.1n 0V)


vA a 0 PWL(0 0V 100n 0V 100.1n 0V 200n 0V 200.1n 0V 300n 0V 300.1n 0V 400n 0V 400.1n 5V
+ 500n 5V 500.1n 5V 600n 5V 600.1n 5V 700n 5V 700.1n 5V 800n 5V 800.1n 0V 900n 0V 900.1n 0V 
+ 1000n 0V 1000.1n 0V 1100n 0V 1100.1n 0V 1200n 0V 1200.1n 5V 1300n 5V 1300.1n 5V 1400n 5V 1400.1n 5V
+ 1500n 5V 1500.1n 5V 1600n 5V 1600.1n 0V 1700n 0V 1700.1n 0V)

VB b 0 PWL(0 0V 100n 0V 100.1n 0V 200n 0V 200.1n 5V 300n 5V 300.1n 5V 400n 5V 400.1n 0V
+ 500n 0V 500.1n 0V 600n 0V 600.1n 5V 700n 5V 700.1n 5V 800n 5V 800.1n 0V 900n 0V 900.1n 0V
+ 1000n 0V 1000.1n 5V 1100n 5V 1100.1n 5V 1200n 5V 1200.1n 0V 1300n 0V 1300.1n 0V 1400n 0V 1400.1n 5V
+ 1500n 5V 1500.1n 5V 1600n 5V 1600.1n 5V 1700n 5V 1700.1n 5V)


***************************************************
* Simulation Options

.options post=2
.tran 1p 1800n


M1000 a_2_100# pin pout Vdd pfet w=9 l=2
+  ad=167 pd=78 as=70 ps=56
M1001 a_2_100# a a_27_101# Vdd pfet w=9 l=2
+  ad=0 pd=0 as=70 ps=56
M1002 a_50_101# abar a_2_100# Vdd pfet w=9 l=2
+  ad=126 pd=46 as=0 ps=0
M1003 vdd b a_50_101# Vdd pfet w=9 l=2
+  ad=426 pd=234 as=0 ps=0
M1004 a_27_101# bbar vdd Vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_18_86# pinbar pout Vdd pfet w=9 l=2
+  ad=161 pd=74 as=0 ps=0
M1006 a_34_86# a a_18_86# Vdd pfet w=9 l=2
+  ad=252 pd=92 as=0 ps=0
M1007 vdd abar a_34_86# Vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_34_86# b vdd Vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_18_86# bbar a_34_86# Vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 pinbar pin vdd Vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 a_50_74# abar vdd Vdd pfet w=8 l=2
+  ad=72 pd=52 as=0 ps=0
M1012 abar a vdd Vdd pfet w=7 l=2
+  ad=29 pd=24 as=0 ps=0
M1013 pinbar pin gnd Gnd nfet w=3 l=2
+  ad=19 pd=18 as=210 ps=172
M1014 a_82_70# bbar vdd Vdd pfet w=8 l=2
+  ad=112 pd=44 as=0 ps=0
M1015 fout min a_82_70# Vdd pfet w=8 l=2
+  ad=112 pd=44 as=0 ps=0
M1016 a_50_74# minbar fout Vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 bbar b vdd Vdd pfet w=7 l=2
+  ad=29 pd=24 as=0 ps=0
M1018 abar a gnd Gnd nfet w=5 l=2
+  ad=23 pd=20 as=0 ps=0
M1019 minbar min vdd Vdd pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1020 bbar b gnd Gnd nfet w=5 l=2
+  ad=23 pd=20 as=0 ps=0
M1021 a_50_31# abar fout Gnd nfet w=4 l=2
+  ad=96 pd=72 as=40 ps=36
M1022 minbar min gnd Gnd nfet w=3 l=2
+  ad=19 pd=18 as=0 ps=0
M1023 gnd bbar a_50_31# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 a_50_31# min gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 fout minbar a_50_31# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 a_2_9# pinbar pout Gnd nfet w=5 l=2
+  ad=162 pd=118 as=93 ps=58
M1027 pout a a_27_23# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=46 ps=40
M1028 a_50_22# abar pout Gnd nfet w=5 l=2
+  ad=70 pd=38 as=0 ps=0
M1029 a_2_9# b a_50_22# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 a_27_23# bbar a_2_9# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 a_2_9# pin gnd Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 a_34_9# a a_2_9# Gnd nfet w=5 l=2
+  ad=140 pd=76 as=0 ps=0
M1033 gnd abar a_34_9# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 a_34_9# b gnd Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 a_2_9# bbar a_34_9# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_2_9# Gnd 2.68fF
C1 a_50_31# Gnd 3.09fF
C2 fout Gnd 6.88fF
C3 minbar Gnd 2.24fF
C4 min Gnd 8.58fF
C5 gnd Gnd 15.60fF
C6 a_50_74# Gnd 2.30fF
C7 pinbar Gnd 2.59fF
C8 bbar Gnd 2.49fF
C9 vdd Gnd 16.34fF
C10 abar Gnd 2.49fF
C11 a_27_101# Gnd 2.09fF
C12 pout Gnd 7.64fF
C13 pin Gnd 3.66fF
