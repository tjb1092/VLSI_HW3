magic
tech scmos
timestamp 1539095088
<< metal1 >>
rect 47 141 51 145
rect 79 141 83 145
rect 186 141 190 145
rect 218 141 222 145
rect 325 141 329 145
rect 357 141 361 145
rect 464 141 468 145
rect 496 141 500 145
rect 603 141 607 145
rect 635 141 639 145
rect 742 141 746 145
rect 774 141 778 145
rect 881 141 885 145
rect 913 141 917 145
rect 1020 141 1024 145
rect 1052 141 1056 145
rect -7 131 0 134
rect 1112 131 1115 134
rect -7 10 -4 131
rect 1112 124 1116 128
rect 1112 13 1116 17
rect -7 7 0 10
rect 1112 7 1115 10
rect 135 -4 139 0
rect 274 -4 278 0
rect 413 -4 417 0
rect 552 -4 556 0
rect 691 -4 695 0
rect 830 -4 834 0
rect 969 -4 973 0
rect 1108 -4 1112 0
use P3_take3  P3_take3_0
array 0 7 139 0 0 141
timestamp 1539012001
transform 1 0 16 0 1 10
box -16 -10 123 131
<< labels >>
rlabel metal1 1112 13 1116 17 7 gnd
rlabel metal1 1112 124 1116 128 7 vdd
rlabel metal1 1112 131 1115 134 7 pin
rlabel metal1 1112 7 1115 10 7 mout
rlabel metal1 1052 141 1056 145 5 b0
rlabel metal1 1020 141 1024 145 5 a0
rlabel metal1 913 141 917 145 5 b1
rlabel metal1 881 141 885 145 5 a1
rlabel metal1 774 141 778 145 5 b2
rlabel metal1 742 141 746 145 5 a2
rlabel metal1 635 141 639 145 5 b3
rlabel metal1 603 141 607 145 5 a3
rlabel metal1 496 141 500 145 5 b4
rlabel metal1 464 141 468 145 5 a4
rlabel metal1 357 141 361 145 5 b5
rlabel metal1 325 141 329 145 5 a5
rlabel metal1 218 141 222 145 5 b6
rlabel metal1 186 141 190 145 5 a6
rlabel metal1 79 141 83 145 5 b7
rlabel metal1 47 141 51 145 5 a7
rlabel metal1 135 -4 139 0 1 c7
rlabel metal1 274 -4 278 0 1 c6
rlabel metal1 413 -4 417 0 1 c5
rlabel metal1 552 -4 556 0 1 c4
rlabel metal1 691 -4 695 0 1 c3
rlabel metal1 830 -4 834 0 1 c2
rlabel metal1 969 -4 973 0 1 c1
rlabel metal1 1108 -4 1112 0 1 c0
<< end >>
